`timescale 1 ns / 100 ps
`include "alu-commands.v"

module testbench();

    reg [3:0] operation = 0;
    reg [31:0] a;
    reg [31:0] b;
    wire [31:0] res;

    alu alu(.a(a), .b(b), .res(res), .operation(operation));
    
    initial begin
        $dumpvars;
        a = 5; b = 3;
        #5 operation = `ALU_NONE;
        #5 operation = `ALU_ADD;
        #5 operation = `ALU_SUB;
        #5 operation = `ALU_XOR;
        #5 operation = `ALU_OR;
        #5 operation = `ALU_AND;
        #5 operation = `ALU_SLL;
        #5 operation = `ALU_SRL;
        #5 operation = `ALU_SRA;
        #5 operation = `ALU_SLT;
        #5 operation = `ALU_SLTU;
        #5 a = 124; b = 45;
        #5 operation = `ALU_NONE;
        #5 operation = `ALU_ADD;
        #5 operation = `ALU_SUB;
        #5 operation = `ALU_XOR;
        #5 operation = `ALU_OR;
        #5 operation = `ALU_AND;
        #5 operation = `ALU_SLL;
        #5 operation = `ALU_SRL;
        #5 operation = `ALU_SRA;
        #5 operation = `ALU_SLT;
        #5 operation = `ALU_SLTU;
        #5 a = 4661; b = 15478;
        #5 operation = `ALU_NONE;
        #5 operation = `ALU_ADD;
        #5 operation = `ALU_SUB;
        #5 operation = `ALU_XOR;
        #5 operation = `ALU_OR;
        #5 operation = `ALU_AND;
        #5 operation = `ALU_SLL;
        #5 operation = `ALU_SRL;
        #5 operation = `ALU_SRA;
        #5 operation = `ALU_SLT;
        #5 operation = `ALU_SLTU;
        #5 a = 4294967295; b = 4294967295;
        #5 operation = `ALU_NONE;
        #5 operation = `ALU_ADD;
        #5 operation = `ALU_SUB;
        #5 operation = `ALU_XOR;
        #5 operation = `ALU_OR;
        #5 operation = `ALU_AND;
        #5 operation = `ALU_SLL;
        #5 operation = `ALU_SRL;
        #5 operation = `ALU_SRA;
        #5 operation = `ALU_SLT;
        #5 operation = `ALU_SLTU;
        #5 a = 4294967295; b = 1;
        #5 operation = `ALU_NONE;
        #5 operation = `ALU_ADD;
        #5 operation = `ALU_SUB;
        #5 operation = `ALU_XOR;
        #5 operation = `ALU_OR;
        #5 operation = `ALU_AND;
        #5 operation = `ALU_SLL;
        #5 operation = `ALU_SRL;
        #5 operation = `ALU_SRA;
        #5 operation = `ALU_SLT;
        #5 operation = `ALU_SLTU;
        #5 a = 4290000000; b = 4294967295;
        #5 operation = `ALU_NONE;
        #5 operation = `ALU_ADD;
        #5 operation = `ALU_SUB;
        #5 operation = `ALU_XOR;
        #5 operation = `ALU_OR;
        #5 operation = `ALU_AND;
        #5 operation = `ALU_SLL;
        #5 operation = `ALU_SRL;
        #5 operation = `ALU_SRA;
        #5 operation = `ALU_SLT;
        #5 operation = `ALU_SLTU;
        #5 a = 4291111111; b = 4290000000;
        #5 operation = `ALU_NONE;
        #5 operation = `ALU_ADD;
        #5 operation = `ALU_SUB;
        #5 operation = `ALU_XOR;
        #5 operation = `ALU_OR;
        #5 operation = `ALU_AND;
        #5 operation = `ALU_SLL;
        #5 operation = `ALU_SRL;
        #5 operation = `ALU_SRA;
        #5 operation = `ALU_SLT;
        #5 operation = `ALU_SLTU;
        #5 a = 429111111; b = 4290000000;
        #5 operation = `ALU_NONE;
        #5 operation = `ALU_ADD;
        #5 operation = `ALU_SUB;
        #5 operation = `ALU_XOR;
        #5 operation = `ALU_OR;
        #5 operation = `ALU_AND;
        #5 operation = `ALU_SLL;
        #5 operation = `ALU_SRL;
        #5 operation = `ALU_SRA;
        #5 operation = `ALU_SLT;
        #5 operation = `ALU_SLTU;
        #5 a = 4291111111; b = 429000000;
        #5 operation = `ALU_NONE;
        #5 operation = `ALU_ADD;
        #5 operation = `ALU_SUB;
        #5 operation = `ALU_XOR;
        #5 operation = `ALU_OR;
        #5 operation = `ALU_AND;
        #5 operation = `ALU_SLL;
        #5 operation = `ALU_SRL;
        #5 operation = `ALU_SRA;
        #5 operation = `ALU_SLT;
        #5 operation = `ALU_SLTU;
        #5; $finish;
    end
    
endmodule
